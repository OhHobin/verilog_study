`timescale 1ns/1ps

module SR_ff();
    
endmodule