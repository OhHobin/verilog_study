`timescale 1ps/1ps

module testbench();

    SR_ff srff(i0, i1, i2, i3, i4, i5, i6, i7, sel, out);
    
endmodule
