`timescale 1ns/1ps

module register();
   
endmodule