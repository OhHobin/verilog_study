`timescale 1ps/1ps

module testbench();

    T_ff Tff();

endmodule
