`timescale 1ns/1ps

module JK_ff();

endmodule