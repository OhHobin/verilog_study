`timescale 1ps/1ps

module testbench();
    

    JK_ff JKff(i0, i1, i2, i3, i4, i5, i6, i7, sel, out);
    
endmodule
