`timescale 1ns/1ps

module T_ff();

endmodule