`timescale 1ps/1ps

module testbench();

    register rreg();
    
endmodule
