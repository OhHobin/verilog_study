`timescale 1ps/1ps

module testbench();

    D_ff Dff();

endmodule
